/*
 Author: Yash Parikh
 File: my_VGA_project_top.v
 Description: Top level module of my DE1-SoC VGA test project
*/

